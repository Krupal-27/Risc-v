`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/04/2025 02:24:45 PM
// Design Name: 
// Module Name: RISC_V
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module pipe_MIPS (clk1, clk2);
 
 input clk1, clk2; // two phase clocks 

 reg [31:0] PC, IF_ID_IR, IF_ID_NPC;
 reg [31:0] ID_EX_IR, ID_EX_NPC, ID_EX_A, ID_EX_B, ID_EX_Imm;
 reg [4:0] ID_EX_type, EX_MEM_type, MEM_WB_type; // INDICATE AND TRASNFER THE INSTRUCTION TYPE
 reg [31:0] EX_MEM_IR, EX_MEM_ALUOut, EX_MEM_B;
 reg EX_MEM_cond;
 reg [31:0] MEM_WB_IR, MEM_WB_ALUOut, MEM_WB_LMD;
 reg [31:0] REG [0:31]; // REGISTER BANK ( 32*32 BITS  )
 reg [31:0] MEM [0:1023]; // data memory

 parameter ADD=6'b000000, SUB=6'b000001, AND=6'b000010, OR=6'b000011, SLT=6'b000100,
           MUL=6'b000101, HLT=6'b111111, LW=6'b001000, SW=6'b001001,
           ADDI=6'b001010, SUBI=6'b001011, ANDI=6'b001100, ORI=6'b001101, SLTI=6'b001110,
           BNEQZ=6'b001111, BEQZ=6'b010000;

parameter RR_ALU=3'b000, RM_ALU=3'b001, LOAD=3'b010, STORE=3'b011, BRANCH=3'b100, HALT=3'b101;

 reg HALTED; // SET AFTER HLT INSTRUCTION IS COMPLETED ( IN WB STAGE)
 reg TAKEN_BRANCH; // SET IF BRANCH IS TAKEN           

 // IF STAGE 
 
 always @(posedge clk1)
   if ( HALTED == 0)
   begin
    if (((EX_MEM_IR[31:26] == BEQZ) && (EX_MEM_cond == 1)) || // WHEN BRANCH IS ACTIVE 
        ((EX_MEM_IR[31:26] == BNEQZ) && (EX_MEM_cond == 0)) )
        begin
            IF_ID_IR <= MEM[EX_MEM_ALUOut];
            TAKEN_BRANCH <= 1'b1;
            IF_ID_NPC <= EX_MEM_ALUOut + 1;
            PC <= EX_MEM_ALUOut + 1;
        end
        else
        begin
            IF_ID_IR <= MEM[PC]; // NORMAL INSTRUCTION FETCH ADD 1
            IF_ID_NPC <= PC + 1;
            PC <= PC + 1;
        end 
   end

   // ID STAGE 

   always @(posedge clk2)
   if ( HALTED == 0)
   begin
    if (IF_ID_IR[25:21] == 5'b00000) ID_EX_A <= 0;
    else ID_EX_A <= REG[IF_ID_IR[25:21]]; // rs stage TAKE FROM REGISTER BANK 

    if (IF_ID_IR[20:16] == 5'b00000) ID_EX_B <= 0;
    else ID_EX_B <= REG[IF_ID_IR[20:16]]; // rt stage TAKE FROM REGISTER BANK

    ID_EX_NPC <= IF_ID_NPC;
    ID_EX_IR <= IF_ID_IR;
    ID_EX_Imm <= {{16{IF_ID_IR[15]}}, IF_ID_IR[15:0]}; // SIGN EXTENSION

    case (IF_ID_IR [31:26])
        ADD, SUB, AND, OR, SLT, MUL: ID_EX_type <= RR_ALU;
        ADDI, SUBI, SLTI           : ID_EX_type <= RM_ALU;
        LW                         : ID_EX_type <= LOAD;
        SW                         : ID_EX_type <= STORE;
        BEQZ, BNEQZ                : ID_EX_type <= BRANCH;
        HLT                        : ID_EX_type <= HALT;
        default                    : ID_EX_type <= HALT; // INVALID OPCODE
    endcase
    end

    // EXECUTION STAGE
     always @ (posedge clk1)
        if ( HALTED == 0)
        begin
            EX_MEM_type <= ID_EX_type;
            EX_MEM_IR <= ID_EX_IR;
            TAKEN_BRANCH <= 0;

            case (ID_EX_type)
                RR_ALU: begin
                            case (ID_EX_IR[31:26])
                                ADD: EX_MEM_ALUOut <= ID_EX_A + ID_EX_B;
                                SUB: EX_MEM_ALUOut <= ID_EX_A - ID_EX_B;
                                AND: EX_MEM_ALUOut <= ID_EX_A & ID_EX_B;
                                OR : EX_MEM_ALUOut <= ID_EX_A | ID_EX_B;
                                SLT: EX_MEM_ALUOut <= ID_EX_A < ID_EX_B;
                                MUL: EX_MEM_ALUOut <= ID_EX_A * ID_EX_B;
                                default: EX_MEM_ALUOut <= 32'hxxxxxxxx; // INVALID OPCODE
                            endcase
                end

                RM_ALU: begin
                            case (ID_EX_IR[31:26]) // OPCODE
                                ADDI: EX_MEM_ALUOut <= ID_EX_A + ID_EX_Imm;
                                SUBI: EX_MEM_ALUOut <= ID_EX_A - ID_EX_Imm;
                                SLTI: EX_MEM_ALUOut <= ID_EX_A < ID_EX_Imm;
                                default: EX_MEM_ALUOut <= 32'hxxxxxxxx; // INVALID OPCODE
                            endcase
                end

                LOAD, STORE: begin
                            EX_MEM_ALUOut <= ID_EX_A + ID_EX_Imm; 
                             EX_MEM_B <= ID_EX_B; // USE FOR NEXT STEP STORE THE VALUE
                end

                BRANCH: begin
                            EX_MEM_ALUOut <= ID_EX_NPC + ID_EX_Imm; 
                            EX_MEM_cond <= (ID_EX_A == 0);
                end
            endcase
        end

// MEMORY STAGE
    always @(posedge clk2)
        if ( HALTED == 0)
        begin
            MEM_WB_type <= EX_MEM_type;
            MEM_WB_IR <= EX_MEM_IR;

            case (EX_MEM_type)
            RR_ALU, RM_ALU: 
                MEM_WB_ALUOut <= EX_MEM_ALUOut;
                
                LOAD: MEM_WB_LMD <= MEM[EX_MEM_ALUOut]; // LOAD THE VALUE FROM MEMORY

                STORE: if (TAKEN_BRANCH == 0) // STORE ONLY IF BRANCH NOT TAKEN
                       MEM[EX_MEM_ALUOut] <= EX_MEM_B;
            endcase
        end

        // WB WRITE BACK STAGE 
        always @(posedge clk1)
        begin
            if (TAKEN_BRANCH == 0) // DISABLE WRITE BACK IF BRANCH TAKEN
            case (MEM_WB_type)
                RR_ALU: REG[MEM_WB_IR[15:11]] <= MEM_WB_ALUOut; // rd field

                RM_ALU: REG[MEM_WB_IR[20:16]] <= MEM_WB_ALUOut; // rt field

                LOAD: REG[MEM_WB_IR[20:16]] <= MEM_WB_LMD; // rt field

                HALT: HALTED <= 1'b1; // SET HALTED FLAG PROCESSOR OFF
            endcase
        end

    
endmodule


